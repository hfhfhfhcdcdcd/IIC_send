module alarm (
    
);
    
endmodule