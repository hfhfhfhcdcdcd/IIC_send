module e2prom_top (
    
);
    
endmodule