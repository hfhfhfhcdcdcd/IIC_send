module  (
    
);
    
endmodule